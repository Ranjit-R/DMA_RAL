  // -------------------------------------------------
  // Global parameters
  // -------------------------------------------------
 `define data_width  32
 `define addr_width  32
