package dma_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  //--------------------------------------------------
  // Sequence_item
  //--------------------------------------------------
  `include "bus_sequence_item.sv"

  // -------------------------------------------------
  // RAL registers
  // -------------------------------------------------
  `include "dma_reg_class.sv"
  `include "top_dma_reg_block.sv"

  // -------------------------------------------------
  // Sequence item & sequencer
  // -------------------------------------------------
  `include "dma_sequence_item.sv"
  `include "dma_sequencer.sv"

  // -------------------------------------------------
  // Driver & Monitor
  // -------------------------------------------------
  `include "dma_driver.sv"
  `include "dma_monitor.sv"

  // -------------------------------------------------
  // Agent
  // -------------------------------------------------
  `include "dma_agent.sv"

  // -------------------------------------------------
  // Scoreboard
  // -------------------------------------------------
  `include "dma_scoreboard.sv"



  // -------------------------------------------------
  // Adapter & sequences
  // -------------------------------------------------
  `include "top_dma_adapter.sv"
  `include "dma_reg_sequence.sv"

  // -------------------------------------------------
  // Environment
  // -------------------------------------------------
  `include "dma_environment.sv"

  // -------------------------------------------------
  // Test
  // -------------------------------------------------
  `include "dma_test.sv"

endpackage : dma_pkg
